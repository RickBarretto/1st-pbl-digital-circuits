module display(
    output top_segment,
    output top_left_segment,
    output top_right_segment,
    output middle_segment,
    output bottom_left_segment,
    output bottom_right_segment,
    output bottom_segment,

    input [2:0] encoded_entry
);


endmodule 