module display(
    output top_segment,
    output top_left_segment,
    output top_right_segment,
    output middle_segment,
    output bottom_left_segment,
    output bottom_right_segment,
    output bottom_segment,

    input irrigation_mode_on,
    
    input conflicting_water_sensor,
    input low_water_level,
    input mid_water_level,
    input high_water_level,

    input dripper, 
    input splinker
);
    

endmodule 